// mityarm_5csx_dev_board_tb.v

// Generated using ACDS version 13.1 162 at 2014.02.17.18:47:33

`timescale 1 ps / 1 ps
module mityarm_5csx_dev_board_tb (
	);

	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_odt;                             // mityarm_5csx_dev_board_inst:hps_ddr_mem_odt -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_odt
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_cs_n;                            // mityarm_5csx_dev_board_inst:hps_ddr_mem_cs_n -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_cs_n
	wire  [14:0] mityarm_5csx_dev_board_inst_hps_ddr_mem_a;                               // mityarm_5csx_dev_board_inst:hps_ddr_mem_a -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_a
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_ddr_bfm_conduit_oct_rzqin;               // mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_oct_rzqin -> mityarm_5csx_dev_board_inst:hps_ddr_oct_rzqin
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_ck_n;                            // mityarm_5csx_dev_board_inst:hps_ddr_mem_ck_n -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_ck_n
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_ras_n;                           // mityarm_5csx_dev_board_inst:hps_ddr_mem_ras_n -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_ras_n
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_cke;                             // mityarm_5csx_dev_board_inst:hps_ddr_mem_cke -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_cke
	wire   [4:0] mityarm_5csx_dev_board_inst_hps_ddr_mem_dqs;                             // [] -> [mityarm_5csx_dev_board_inst:hps_ddr_mem_dqs, mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_dqs]
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_we_n;                            // mityarm_5csx_dev_board_inst:hps_ddr_mem_we_n -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_we_n
	wire   [2:0] mityarm_5csx_dev_board_inst_hps_ddr_mem_ba;                              // mityarm_5csx_dev_board_inst:hps_ddr_mem_ba -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_ba
	wire  [39:0] mityarm_5csx_dev_board_inst_hps_ddr_mem_dq;                              // [] -> [mityarm_5csx_dev_board_inst:hps_ddr_mem_dq, mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_dq]
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_ck;                              // mityarm_5csx_dev_board_inst:hps_ddr_mem_ck -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_ck
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_reset_n;                         // mityarm_5csx_dev_board_inst:hps_ddr_mem_reset_n -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_reset_n
	wire   [4:0] mityarm_5csx_dev_board_inst_hps_ddr_mem_dm;                              // mityarm_5csx_dev_board_inst:hps_ddr_mem_dm -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_dm
	wire         mityarm_5csx_dev_board_inst_hps_ddr_mem_cas_n;                           // mityarm_5csx_dev_board_inst:hps_ddr_mem_cas_n -> mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_cas_n
	wire   [4:0] mityarm_5csx_dev_board_inst_hps_ddr_mem_dqs_n;                           // [] -> [mityarm_5csx_dev_board_inst:hps_ddr_mem_dqs_n, mityarm_5csx_dev_board_inst_hps_ddr_bfm:sig_mem_dqs_n]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c0_inst_sda;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_i2c0_inst_SDA, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_i2c0_inst_SDA]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_tx_ctl;             // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_TX_CTL -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_TX_CTL
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_mdio;               // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_MDIO, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_MDIO]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio28;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO28, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO28]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c0_inst_scl;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_i2c0_inst_SCL, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_i2c0_inst_SCL]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d5;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D5, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D5]
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_clk;     // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_CLK -> mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_CLK
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d4;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D4, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D4]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d7;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D7, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D7]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d6;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D6, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D6]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d1;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D1, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D1]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_can1_inst_tx;                  // mityarm_5csx_dev_board_inst:hps_io_hps_io_can1_inst_TX -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_can1_inst_TX
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d0;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D0, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D0]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d3;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D3, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D3]
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rx_clk; // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_RX_CLK -> mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_RX_CLK
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d2;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_D2, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_D2]
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_can0_inst_rx;      // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_can0_inst_RX -> mityarm_5csx_dev_board_inst:hps_io_hps_io_can0_inst_RX
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_uart0_inst_rx;     // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_uart0_inst_RX -> mityarm_5csx_dev_board_inst:hps_io_hps_io_uart0_inst_RX
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd3;   // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_RXD3 -> mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_RXD3
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd2;   // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_RXD2 -> mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_RXD2
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c1_inst_scl;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_i2c1_inst_SCL, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_i2c1_inst_SCL]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio50;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO50, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO50]
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rx_ctl; // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_RX_CTL -> mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_RX_CTL
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_stp;                 // mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_STP -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_STP
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_clk;                 // mityarm_5csx_dev_board_inst:hps_io_hps_io_sdio_inst_CLK -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_sdio_inst_CLK
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d1;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_sdio_inst_D1, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_sdio_inst_D1]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d0;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_sdio_inst_D0, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_sdio_inst_D0]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d3;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_sdio_inst_D3, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_sdio_inst_D3]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d2;                  // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_sdio_inst_D2, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_sdio_inst_D2]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio48;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO48, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO48]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio00;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO00, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO00]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio49;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO49, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO49]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io3;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_IO3, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_IO3]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd1;               // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_TXD1 -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_TXD1
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io2;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_IO2, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_IO2]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd0;               // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_TXD0 -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_TXD0
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io1;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_IO1, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_IO1]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd3;               // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_TXD3 -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_TXD3
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io0;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_IO0, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_IO0]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd2;               // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_TXD2 -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_TXD2
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_dir;     // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_DIR -> mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_DIR
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd0;   // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_RXD0 -> mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_RXD0
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c1_inst_sda;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_i2c1_inst_SDA, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_i2c1_inst_SDA]
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd1;   // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_RXD1 -> mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_RXD1
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_cmd;                 // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_sdio_inst_CMD, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_sdio_inst_CMD]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_clk;                 // mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_CLK -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_CLK
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio41;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO41, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO41]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio09;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO09, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO09]
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_can1_inst_rx;      // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_can1_inst_RX -> mityarm_5csx_dev_board_inst:hps_io_hps_io_can1_inst_RX
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio40;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO40, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO40]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_mdc;                // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_MDC -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_MDC
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio37;              // [] -> [mityarm_5csx_dev_board_inst:hps_io_hps_io_gpio_inst_GPIO37, mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_gpio_inst_GPIO37]
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_uart0_inst_tx;                 // mityarm_5csx_dev_board_inst:hps_io_hps_io_uart0_inst_TX -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_uart0_inst_TX
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_can0_inst_tx;                  // mityarm_5csx_dev_board_inst:hps_io_hps_io_can0_inst_TX -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_can0_inst_TX
	wire   [0:0] mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_nxt;     // mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_usb1_inst_NXT -> mityarm_5csx_dev_board_inst:hps_io_hps_io_usb1_inst_NXT
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_ss1;                 // mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_SS1 -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_SS1
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_tx_clk;             // mityarm_5csx_dev_board_inst:hps_io_hps_io_emac1_inst_TX_CLK -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_emac1_inst_TX_CLK
	wire         mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_ss0;                 // mityarm_5csx_dev_board_inst:hps_io_hps_io_qspi_inst_SS0 -> mityarm_5csx_dev_board_inst_hps_io_bfm:sig_hps_io_qspi_inst_SS0

	mityarm_5csx_dev_board mityarm_5csx_dev_board_inst (
		.hps_ddr_mem_a                   (mityarm_5csx_dev_board_inst_hps_ddr_mem_a),                               // hps_ddr.mem_a
		.hps_ddr_mem_ba                  (mityarm_5csx_dev_board_inst_hps_ddr_mem_ba),                              //        .mem_ba
		.hps_ddr_mem_ck                  (mityarm_5csx_dev_board_inst_hps_ddr_mem_ck),                              //        .mem_ck
		.hps_ddr_mem_ck_n                (mityarm_5csx_dev_board_inst_hps_ddr_mem_ck_n),                            //        .mem_ck_n
		.hps_ddr_mem_cke                 (mityarm_5csx_dev_board_inst_hps_ddr_mem_cke),                             //        .mem_cke
		.hps_ddr_mem_cs_n                (mityarm_5csx_dev_board_inst_hps_ddr_mem_cs_n),                            //        .mem_cs_n
		.hps_ddr_mem_ras_n               (mityarm_5csx_dev_board_inst_hps_ddr_mem_ras_n),                           //        .mem_ras_n
		.hps_ddr_mem_cas_n               (mityarm_5csx_dev_board_inst_hps_ddr_mem_cas_n),                           //        .mem_cas_n
		.hps_ddr_mem_we_n                (mityarm_5csx_dev_board_inst_hps_ddr_mem_we_n),                            //        .mem_we_n
		.hps_ddr_mem_reset_n             (mityarm_5csx_dev_board_inst_hps_ddr_mem_reset_n),                         //        .mem_reset_n
		.hps_ddr_mem_dq                  (mityarm_5csx_dev_board_inst_hps_ddr_mem_dq),                              //        .mem_dq
		.hps_ddr_mem_dqs                 (mityarm_5csx_dev_board_inst_hps_ddr_mem_dqs),                             //        .mem_dqs
		.hps_ddr_mem_dqs_n               (mityarm_5csx_dev_board_inst_hps_ddr_mem_dqs_n),                           //        .mem_dqs_n
		.hps_ddr_mem_odt                 (mityarm_5csx_dev_board_inst_hps_ddr_mem_odt),                             //        .mem_odt
		.hps_ddr_mem_dm                  (mityarm_5csx_dev_board_inst_hps_ddr_mem_dm),                              //        .mem_dm
		.hps_ddr_oct_rzqin               (mityarm_5csx_dev_board_inst_hps_ddr_bfm_conduit_oct_rzqin),               //        .oct_rzqin
		.hps_io_hps_io_emac1_inst_TX_CLK (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_tx_clk),             //  hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_hps_io_emac1_inst_TXD0   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd0),               //        .hps_io_emac1_inst_TXD0
		.hps_io_hps_io_emac1_inst_TXD1   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd1),               //        .hps_io_emac1_inst_TXD1
		.hps_io_hps_io_emac1_inst_TXD2   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd2),               //        .hps_io_emac1_inst_TXD2
		.hps_io_hps_io_emac1_inst_TXD3   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd3),               //        .hps_io_emac1_inst_TXD3
		.hps_io_hps_io_emac1_inst_RXD0   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd0),   //        .hps_io_emac1_inst_RXD0
		.hps_io_hps_io_emac1_inst_MDIO   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_mdio),               //        .hps_io_emac1_inst_MDIO
		.hps_io_hps_io_emac1_inst_MDC    (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_mdc),                //        .hps_io_emac1_inst_MDC
		.hps_io_hps_io_emac1_inst_RX_CTL (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rx_ctl), //        .hps_io_emac1_inst_RX_CTL
		.hps_io_hps_io_emac1_inst_TX_CTL (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_tx_ctl),             //        .hps_io_emac1_inst_TX_CTL
		.hps_io_hps_io_emac1_inst_RX_CLK (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rx_clk), //        .hps_io_emac1_inst_RX_CLK
		.hps_io_hps_io_emac1_inst_RXD1   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd1),   //        .hps_io_emac1_inst_RXD1
		.hps_io_hps_io_emac1_inst_RXD2   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd2),   //        .hps_io_emac1_inst_RXD2
		.hps_io_hps_io_emac1_inst_RXD3   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd3),   //        .hps_io_emac1_inst_RXD3
		.hps_io_hps_io_qspi_inst_SS1     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_ss1),                 //        .hps_io_qspi_inst_SS1
		.hps_io_hps_io_qspi_inst_IO0     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io0),                 //        .hps_io_qspi_inst_IO0
		.hps_io_hps_io_qspi_inst_IO1     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io1),                 //        .hps_io_qspi_inst_IO1
		.hps_io_hps_io_qspi_inst_IO2     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io2),                 //        .hps_io_qspi_inst_IO2
		.hps_io_hps_io_qspi_inst_IO3     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io3),                 //        .hps_io_qspi_inst_IO3
		.hps_io_hps_io_qspi_inst_SS0     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_ss0),                 //        .hps_io_qspi_inst_SS0
		.hps_io_hps_io_qspi_inst_CLK     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_clk),                 //        .hps_io_qspi_inst_CLK
		.hps_io_hps_io_sdio_inst_CMD     (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_cmd),                 //        .hps_io_sdio_inst_CMD
		.hps_io_hps_io_sdio_inst_D0      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d0),                  //        .hps_io_sdio_inst_D0
		.hps_io_hps_io_sdio_inst_D1      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d1),                  //        .hps_io_sdio_inst_D1
		.hps_io_hps_io_sdio_inst_CLK     (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_clk),                 //        .hps_io_sdio_inst_CLK
		.hps_io_hps_io_sdio_inst_D2      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d2),                  //        .hps_io_sdio_inst_D2
		.hps_io_hps_io_sdio_inst_D3      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d3),                  //        .hps_io_sdio_inst_D3
		.hps_io_hps_io_usb1_inst_D0      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d0),                  //        .hps_io_usb1_inst_D0
		.hps_io_hps_io_usb1_inst_D1      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d1),                  //        .hps_io_usb1_inst_D1
		.hps_io_hps_io_usb1_inst_D2      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d2),                  //        .hps_io_usb1_inst_D2
		.hps_io_hps_io_usb1_inst_D3      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d3),                  //        .hps_io_usb1_inst_D3
		.hps_io_hps_io_usb1_inst_D4      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d4),                  //        .hps_io_usb1_inst_D4
		.hps_io_hps_io_usb1_inst_D5      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d5),                  //        .hps_io_usb1_inst_D5
		.hps_io_hps_io_usb1_inst_D6      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d6),                  //        .hps_io_usb1_inst_D6
		.hps_io_hps_io_usb1_inst_D7      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d7),                  //        .hps_io_usb1_inst_D7
		.hps_io_hps_io_usb1_inst_CLK     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_clk),     //        .hps_io_usb1_inst_CLK
		.hps_io_hps_io_usb1_inst_STP     (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_stp),                 //        .hps_io_usb1_inst_STP
		.hps_io_hps_io_usb1_inst_DIR     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_dir),     //        .hps_io_usb1_inst_DIR
		.hps_io_hps_io_usb1_inst_NXT     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_nxt),     //        .hps_io_usb1_inst_NXT
		.hps_io_hps_io_uart0_inst_RX     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_uart0_inst_rx),     //        .hps_io_uart0_inst_RX
		.hps_io_hps_io_uart0_inst_TX     (mityarm_5csx_dev_board_inst_hps_io_hps_io_uart0_inst_tx),                 //        .hps_io_uart0_inst_TX
		.hps_io_hps_io_i2c0_inst_SDA     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c0_inst_sda),                 //        .hps_io_i2c0_inst_SDA
		.hps_io_hps_io_i2c0_inst_SCL     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c0_inst_scl),                 //        .hps_io_i2c0_inst_SCL
		.hps_io_hps_io_i2c1_inst_SDA     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c1_inst_sda),                 //        .hps_io_i2c1_inst_SDA
		.hps_io_hps_io_i2c1_inst_SCL     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c1_inst_scl),                 //        .hps_io_i2c1_inst_SCL
		.hps_io_hps_io_can0_inst_RX      (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_can0_inst_rx),      //        .hps_io_can0_inst_RX
		.hps_io_hps_io_can0_inst_TX      (mityarm_5csx_dev_board_inst_hps_io_hps_io_can0_inst_tx),                  //        .hps_io_can0_inst_TX
		.hps_io_hps_io_can1_inst_RX      (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_can1_inst_rx),      //        .hps_io_can1_inst_RX
		.hps_io_hps_io_can1_inst_TX      (mityarm_5csx_dev_board_inst_hps_io_hps_io_can1_inst_tx),                  //        .hps_io_can1_inst_TX
		.hps_io_hps_io_gpio_inst_GPIO00  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio00),              //        .hps_io_gpio_inst_GPIO00
		.hps_io_hps_io_gpio_inst_GPIO09  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio09),              //        .hps_io_gpio_inst_GPIO09
		.hps_io_hps_io_gpio_inst_GPIO28  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio28),              //        .hps_io_gpio_inst_GPIO28
		.hps_io_hps_io_gpio_inst_GPIO37  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio37),              //        .hps_io_gpio_inst_GPIO37
		.hps_io_hps_io_gpio_inst_GPIO40  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio40),              //        .hps_io_gpio_inst_GPIO40
		.hps_io_hps_io_gpio_inst_GPIO41  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio41),              //        .hps_io_gpio_inst_GPIO41
		.hps_io_hps_io_gpio_inst_GPIO48  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio48),              //        .hps_io_gpio_inst_GPIO48
		.hps_io_hps_io_gpio_inst_GPIO49  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio49),              //        .hps_io_gpio_inst_GPIO49
		.hps_io_hps_io_gpio_inst_GPIO50  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio50)               //        .hps_io_gpio_inst_GPIO50
	);

	altera_conduit_bfm mityarm_5csx_dev_board_inst_hps_ddr_bfm (
		.sig_mem_a       (mityarm_5csx_dev_board_inst_hps_ddr_mem_a),                 // conduit.mem_a
		.sig_mem_ba      (mityarm_5csx_dev_board_inst_hps_ddr_mem_ba),                //        .mem_ba
		.sig_mem_ck      (mityarm_5csx_dev_board_inst_hps_ddr_mem_ck),                //        .mem_ck
		.sig_mem_ck_n    (mityarm_5csx_dev_board_inst_hps_ddr_mem_ck_n),              //        .mem_ck_n
		.sig_mem_cke     (mityarm_5csx_dev_board_inst_hps_ddr_mem_cke),               //        .mem_cke
		.sig_mem_cs_n    (mityarm_5csx_dev_board_inst_hps_ddr_mem_cs_n),              //        .mem_cs_n
		.sig_mem_ras_n   (mityarm_5csx_dev_board_inst_hps_ddr_mem_ras_n),             //        .mem_ras_n
		.sig_mem_cas_n   (mityarm_5csx_dev_board_inst_hps_ddr_mem_cas_n),             //        .mem_cas_n
		.sig_mem_we_n    (mityarm_5csx_dev_board_inst_hps_ddr_mem_we_n),              //        .mem_we_n
		.sig_mem_reset_n (mityarm_5csx_dev_board_inst_hps_ddr_mem_reset_n),           //        .mem_reset_n
		.sig_mem_dq      (mityarm_5csx_dev_board_inst_hps_ddr_mem_dq),                //        .mem_dq
		.sig_mem_dqs     (mityarm_5csx_dev_board_inst_hps_ddr_mem_dqs),               //        .mem_dqs
		.sig_mem_dqs_n   (mityarm_5csx_dev_board_inst_hps_ddr_mem_dqs_n),             //        .mem_dqs_n
		.sig_mem_odt     (mityarm_5csx_dev_board_inst_hps_ddr_mem_odt),               //        .mem_odt
		.sig_mem_dm      (mityarm_5csx_dev_board_inst_hps_ddr_mem_dm),                //        .mem_dm
		.sig_oct_rzqin   (mityarm_5csx_dev_board_inst_hps_ddr_bfm_conduit_oct_rzqin)  //        .oct_rzqin
	);

	altera_conduit_bfm_0002 mityarm_5csx_dev_board_inst_hps_io_bfm (
		.sig_hps_io_emac1_inst_TX_CLK (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_tx_clk),             // conduit.hps_io_emac1_inst_TX_CLK
		.sig_hps_io_emac1_inst_TXD0   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd0),               //        .hps_io_emac1_inst_TXD0
		.sig_hps_io_emac1_inst_TXD1   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd1),               //        .hps_io_emac1_inst_TXD1
		.sig_hps_io_emac1_inst_TXD2   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd2),               //        .hps_io_emac1_inst_TXD2
		.sig_hps_io_emac1_inst_TXD3   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_txd3),               //        .hps_io_emac1_inst_TXD3
		.sig_hps_io_emac1_inst_RXD0   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd0),   //        .hps_io_emac1_inst_RXD0
		.sig_hps_io_emac1_inst_MDIO   (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_mdio),               //        .hps_io_emac1_inst_MDIO
		.sig_hps_io_emac1_inst_MDC    (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_mdc),                //        .hps_io_emac1_inst_MDC
		.sig_hps_io_emac1_inst_RX_CTL (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rx_ctl), //        .hps_io_emac1_inst_RX_CTL
		.sig_hps_io_emac1_inst_TX_CTL (mityarm_5csx_dev_board_inst_hps_io_hps_io_emac1_inst_tx_ctl),             //        .hps_io_emac1_inst_TX_CTL
		.sig_hps_io_emac1_inst_RX_CLK (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rx_clk), //        .hps_io_emac1_inst_RX_CLK
		.sig_hps_io_emac1_inst_RXD1   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd1),   //        .hps_io_emac1_inst_RXD1
		.sig_hps_io_emac1_inst_RXD2   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd2),   //        .hps_io_emac1_inst_RXD2
		.sig_hps_io_emac1_inst_RXD3   (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_emac1_inst_rxd3),   //        .hps_io_emac1_inst_RXD3
		.sig_hps_io_qspi_inst_SS1     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_ss1),                 //        .hps_io_qspi_inst_SS1
		.sig_hps_io_qspi_inst_IO0     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io0),                 //        .hps_io_qspi_inst_IO0
		.sig_hps_io_qspi_inst_IO1     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io1),                 //        .hps_io_qspi_inst_IO1
		.sig_hps_io_qspi_inst_IO2     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io2),                 //        .hps_io_qspi_inst_IO2
		.sig_hps_io_qspi_inst_IO3     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_io3),                 //        .hps_io_qspi_inst_IO3
		.sig_hps_io_qspi_inst_SS0     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_ss0),                 //        .hps_io_qspi_inst_SS0
		.sig_hps_io_qspi_inst_CLK     (mityarm_5csx_dev_board_inst_hps_io_hps_io_qspi_inst_clk),                 //        .hps_io_qspi_inst_CLK
		.sig_hps_io_sdio_inst_CMD     (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_cmd),                 //        .hps_io_sdio_inst_CMD
		.sig_hps_io_sdio_inst_D0      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d0),                  //        .hps_io_sdio_inst_D0
		.sig_hps_io_sdio_inst_D1      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d1),                  //        .hps_io_sdio_inst_D1
		.sig_hps_io_sdio_inst_CLK     (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_clk),                 //        .hps_io_sdio_inst_CLK
		.sig_hps_io_sdio_inst_D2      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d2),                  //        .hps_io_sdio_inst_D2
		.sig_hps_io_sdio_inst_D3      (mityarm_5csx_dev_board_inst_hps_io_hps_io_sdio_inst_d3),                  //        .hps_io_sdio_inst_D3
		.sig_hps_io_usb1_inst_D0      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d0),                  //        .hps_io_usb1_inst_D0
		.sig_hps_io_usb1_inst_D1      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d1),                  //        .hps_io_usb1_inst_D1
		.sig_hps_io_usb1_inst_D2      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d2),                  //        .hps_io_usb1_inst_D2
		.sig_hps_io_usb1_inst_D3      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d3),                  //        .hps_io_usb1_inst_D3
		.sig_hps_io_usb1_inst_D4      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d4),                  //        .hps_io_usb1_inst_D4
		.sig_hps_io_usb1_inst_D5      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d5),                  //        .hps_io_usb1_inst_D5
		.sig_hps_io_usb1_inst_D6      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d6),                  //        .hps_io_usb1_inst_D6
		.sig_hps_io_usb1_inst_D7      (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_d7),                  //        .hps_io_usb1_inst_D7
		.sig_hps_io_usb1_inst_CLK     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_clk),     //        .hps_io_usb1_inst_CLK
		.sig_hps_io_usb1_inst_STP     (mityarm_5csx_dev_board_inst_hps_io_hps_io_usb1_inst_stp),                 //        .hps_io_usb1_inst_STP
		.sig_hps_io_usb1_inst_DIR     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_dir),     //        .hps_io_usb1_inst_DIR
		.sig_hps_io_usb1_inst_NXT     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_usb1_inst_nxt),     //        .hps_io_usb1_inst_NXT
		.sig_hps_io_uart0_inst_RX     (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_uart0_inst_rx),     //        .hps_io_uart0_inst_RX
		.sig_hps_io_uart0_inst_TX     (mityarm_5csx_dev_board_inst_hps_io_hps_io_uart0_inst_tx),                 //        .hps_io_uart0_inst_TX
		.sig_hps_io_i2c0_inst_SDA     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c0_inst_sda),                 //        .hps_io_i2c0_inst_SDA
		.sig_hps_io_i2c0_inst_SCL     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c0_inst_scl),                 //        .hps_io_i2c0_inst_SCL
		.sig_hps_io_i2c1_inst_SDA     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c1_inst_sda),                 //        .hps_io_i2c1_inst_SDA
		.sig_hps_io_i2c1_inst_SCL     (mityarm_5csx_dev_board_inst_hps_io_hps_io_i2c1_inst_scl),                 //        .hps_io_i2c1_inst_SCL
		.sig_hps_io_can0_inst_RX      (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_can0_inst_rx),      //        .hps_io_can0_inst_RX
		.sig_hps_io_can0_inst_TX      (mityarm_5csx_dev_board_inst_hps_io_hps_io_can0_inst_tx),                  //        .hps_io_can0_inst_TX
		.sig_hps_io_can1_inst_RX      (mityarm_5csx_dev_board_inst_hps_io_bfm_conduit_hps_io_can1_inst_rx),      //        .hps_io_can1_inst_RX
		.sig_hps_io_can1_inst_TX      (mityarm_5csx_dev_board_inst_hps_io_hps_io_can1_inst_tx),                  //        .hps_io_can1_inst_TX
		.sig_hps_io_gpio_inst_GPIO00  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio00),              //        .hps_io_gpio_inst_GPIO00
		.sig_hps_io_gpio_inst_GPIO09  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio09),              //        .hps_io_gpio_inst_GPIO09
		.sig_hps_io_gpio_inst_GPIO28  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio28),              //        .hps_io_gpio_inst_GPIO28
		.sig_hps_io_gpio_inst_GPIO37  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio37),              //        .hps_io_gpio_inst_GPIO37
		.sig_hps_io_gpio_inst_GPIO40  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio40),              //        .hps_io_gpio_inst_GPIO40
		.sig_hps_io_gpio_inst_GPIO41  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio41),              //        .hps_io_gpio_inst_GPIO41
		.sig_hps_io_gpio_inst_GPIO48  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio48),              //        .hps_io_gpio_inst_GPIO48
		.sig_hps_io_gpio_inst_GPIO49  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio49),              //        .hps_io_gpio_inst_GPIO49
		.sig_hps_io_gpio_inst_GPIO50  (mityarm_5csx_dev_board_inst_hps_io_hps_io_gpio_inst_gpio50)               //        .hps_io_gpio_inst_GPIO50
	);

endmodule
