// st_bfm_qsys_tutorial_tb.v

// Generated using ACDS version 13.1 162 at 2014.02.18.10:24:13

`timescale 1 ps / 1 ps
module st_bfm_qsys_tutorial_tb (
	);

	wire         st_bfm_qsys_tutorial_inst_clk_bfm_clk_clk;             // st_bfm_qsys_tutorial_inst_clk_bfm:clk -> [st_bfm_qsys_tutorial_inst:clk_clk, st_bfm_qsys_tutorial_inst_reset_bfm:clk, st_bfm_qsys_tutorial_inst_st_in_bfm:clk, st_bfm_qsys_tutorial_inst_st_out_bfm:clk]
	wire         st_bfm_qsys_tutorial_inst_reset_bfm_reset_reset;       // st_bfm_qsys_tutorial_inst_reset_bfm:reset -> [st_bfm_qsys_tutorial_inst:reset_reset, st_bfm_qsys_tutorial_inst_st_in_bfm:reset, st_bfm_qsys_tutorial_inst_st_out_bfm:reset]
	wire   [0:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_endofpacket;   // st_bfm_qsys_tutorial_inst_st_in_bfm:src_endofpacket -> st_bfm_qsys_tutorial_inst:st_in_endofpacket
	wire   [0:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_valid;         // st_bfm_qsys_tutorial_inst_st_in_bfm:src_valid -> st_bfm_qsys_tutorial_inst:st_in_valid
	wire   [0:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_startofpacket; // st_bfm_qsys_tutorial_inst_st_in_bfm:src_startofpacket -> st_bfm_qsys_tutorial_inst:st_in_startofpacket
	wire   [2:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_error;         // st_bfm_qsys_tutorial_inst_st_in_bfm:src_error -> st_bfm_qsys_tutorial_inst:st_in_error
	wire   [1:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_empty;         // st_bfm_qsys_tutorial_inst_st_in_bfm:src_empty -> st_bfm_qsys_tutorial_inst:st_in_empty
	wire  [31:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_data;          // st_bfm_qsys_tutorial_inst_st_in_bfm:src_data -> st_bfm_qsys_tutorial_inst:st_in_data
	wire   [2:0] st_bfm_qsys_tutorial_inst_st_in_bfm_src_channel;       // st_bfm_qsys_tutorial_inst_st_in_bfm:src_channel -> st_bfm_qsys_tutorial_inst:st_in_channel
	wire         st_bfm_qsys_tutorial_inst_st_in_bfm_src_ready;         // st_bfm_qsys_tutorial_inst:st_in_ready -> st_bfm_qsys_tutorial_inst_st_in_bfm:src_ready
	wire         st_bfm_qsys_tutorial_inst_st_out_endofpacket;          // st_bfm_qsys_tutorial_inst:st_out_endofpacket -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_endofpacket
	wire         st_bfm_qsys_tutorial_inst_st_out_valid;                // st_bfm_qsys_tutorial_inst:st_out_valid -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_valid
	wire         st_bfm_qsys_tutorial_inst_st_out_startofpacket;        // st_bfm_qsys_tutorial_inst:st_out_startofpacket -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_startofpacket
	wire   [2:0] st_bfm_qsys_tutorial_inst_st_out_error;                // st_bfm_qsys_tutorial_inst:st_out_error -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_error
	wire   [1:0] st_bfm_qsys_tutorial_inst_st_out_empty;                // st_bfm_qsys_tutorial_inst:st_out_empty -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_empty
	wire  [31:0] st_bfm_qsys_tutorial_inst_st_out_data;                 // st_bfm_qsys_tutorial_inst:st_out_data -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_data
	wire   [2:0] st_bfm_qsys_tutorial_inst_st_out_channel;              // st_bfm_qsys_tutorial_inst:st_out_channel -> st_bfm_qsys_tutorial_inst_st_out_bfm:sink_channel
	wire         st_bfm_qsys_tutorial_inst_st_out_ready;                // st_bfm_qsys_tutorial_inst_st_out_bfm:sink_ready -> st_bfm_qsys_tutorial_inst:st_out_ready

	st_bfm_qsys_tutorial st_bfm_qsys_tutorial_inst (
		.clk_clk              (st_bfm_qsys_tutorial_inst_clk_bfm_clk_clk),             //    clk.clk
		.reset_reset          (st_bfm_qsys_tutorial_inst_reset_bfm_reset_reset),       //  reset.reset
		.st_in_data           (st_bfm_qsys_tutorial_inst_st_in_bfm_src_data),          //  st_in.data
		.st_in_valid          (st_bfm_qsys_tutorial_inst_st_in_bfm_src_valid),         //       .valid
		.st_in_ready          (st_bfm_qsys_tutorial_inst_st_in_bfm_src_ready),         //       .ready
		.st_in_startofpacket  (st_bfm_qsys_tutorial_inst_st_in_bfm_src_startofpacket), //       .startofpacket
		.st_in_endofpacket    (st_bfm_qsys_tutorial_inst_st_in_bfm_src_endofpacket),   //       .endofpacket
		.st_in_empty          (st_bfm_qsys_tutorial_inst_st_in_bfm_src_empty),         //       .empty
		.st_in_error          (st_bfm_qsys_tutorial_inst_st_in_bfm_src_error),         //       .error
		.st_in_channel        (st_bfm_qsys_tutorial_inst_st_in_bfm_src_channel),       //       .channel
		.st_out_data          (st_bfm_qsys_tutorial_inst_st_out_data),                 // st_out.data
		.st_out_valid         (st_bfm_qsys_tutorial_inst_st_out_valid),                //       .valid
		.st_out_ready         (st_bfm_qsys_tutorial_inst_st_out_ready),                //       .ready
		.st_out_startofpacket (st_bfm_qsys_tutorial_inst_st_out_startofpacket),        //       .startofpacket
		.st_out_endofpacket   (st_bfm_qsys_tutorial_inst_st_out_endofpacket),          //       .endofpacket
		.st_out_empty         (st_bfm_qsys_tutorial_inst_st_out_empty),                //       .empty
		.st_out_error         (st_bfm_qsys_tutorial_inst_st_out_error),                //       .error
		.st_out_channel       (st_bfm_qsys_tutorial_inst_st_out_channel)               //       .channel
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) st_bfm_qsys_tutorial_inst_clk_bfm (
		.clk (st_bfm_qsys_tutorial_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (1),
		.INITIAL_RESET_CYCLES (50)
	) st_bfm_qsys_tutorial_inst_reset_bfm (
		.reset (st_bfm_qsys_tutorial_inst_reset_bfm_reset_reset), // reset.reset
		.clk   (st_bfm_qsys_tutorial_inst_clk_bfm_clk_clk)        //   clk.clk
	);

	altera_avalon_st_source_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (1),
		.USE_ERROR        (1),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (3),
		.ST_ERROR_W       (3),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (7),
		.VHDL_ID          (0)
	) st_bfm_qsys_tutorial_inst_st_in_bfm (
		.clk               (st_bfm_qsys_tutorial_inst_clk_bfm_clk_clk),             //       clk.clk
		.reset             (st_bfm_qsys_tutorial_inst_reset_bfm_reset_reset),       // clk_reset.reset
		.src_data          (st_bfm_qsys_tutorial_inst_st_in_bfm_src_data),          //       src.data
		.src_valid         (st_bfm_qsys_tutorial_inst_st_in_bfm_src_valid),         //          .valid
		.src_ready         (st_bfm_qsys_tutorial_inst_st_in_bfm_src_ready),         //          .ready
		.src_startofpacket (st_bfm_qsys_tutorial_inst_st_in_bfm_src_startofpacket), //          .startofpacket
		.src_endofpacket   (st_bfm_qsys_tutorial_inst_st_in_bfm_src_endofpacket),   //          .endofpacket
		.src_empty         (st_bfm_qsys_tutorial_inst_st_in_bfm_src_empty),         //          .empty
		.src_channel       (st_bfm_qsys_tutorial_inst_st_in_bfm_src_channel),       //          .channel
		.src_error         (st_bfm_qsys_tutorial_inst_st_in_bfm_src_error)          //          .error
	);

	altera_avalon_st_sink_bfm #(
		.USE_PACKET       (1),
		.USE_CHANNEL      (1),
		.USE_ERROR        (1),
		.USE_READY        (1),
		.USE_VALID        (1),
		.USE_EMPTY        (1),
		.ST_SYMBOL_W      (8),
		.ST_NUMSYMBOLS    (4),
		.ST_CHANNEL_W     (3),
		.ST_ERROR_W       (3),
		.ST_EMPTY_W       (2),
		.ST_READY_LATENCY (0),
		.ST_BEATSPERCYCLE (1),
		.ST_MAX_CHANNELS  (7),
		.VHDL_ID          (0)
	) st_bfm_qsys_tutorial_inst_st_out_bfm (
		.clk                (st_bfm_qsys_tutorial_inst_clk_bfm_clk_clk),       //       clk.clk
		.reset              (st_bfm_qsys_tutorial_inst_reset_bfm_reset_reset), // clk_reset.reset
		.sink_data          (st_bfm_qsys_tutorial_inst_st_out_data),           //      sink.data
		.sink_valid         (st_bfm_qsys_tutorial_inst_st_out_valid),          //          .valid
		.sink_ready         (st_bfm_qsys_tutorial_inst_st_out_ready),          //          .ready
		.sink_startofpacket (st_bfm_qsys_tutorial_inst_st_out_startofpacket),  //          .startofpacket
		.sink_endofpacket   (st_bfm_qsys_tutorial_inst_st_out_endofpacket),    //          .endofpacket
		.sink_empty         (st_bfm_qsys_tutorial_inst_st_out_empty),          //          .empty
		.sink_channel       (st_bfm_qsys_tutorial_inst_st_out_channel),        //          .channel
		.sink_error         (st_bfm_qsys_tutorial_inst_st_out_error)           //          .error
	);

endmodule
