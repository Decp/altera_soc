// st_bfm_qsys_tutorial.v

// Generated using ACDS version 13.1 162 at 2014.02.18.10:24:14

`timescale 1 ps / 1 ps
module st_bfm_qsys_tutorial (
		input  wire        clk_clk,              //    clk.clk
		input  wire        reset_reset,          //  reset.reset
		input  wire [31:0] st_in_data,           //  st_in.data
		input  wire        st_in_valid,          //       .valid
		output wire        st_in_ready,          //       .ready
		input  wire        st_in_startofpacket,  //       .startofpacket
		input  wire        st_in_endofpacket,    //       .endofpacket
		input  wire [1:0]  st_in_empty,          //       .empty
		input  wire [2:0]  st_in_error,          //       .error
		input  wire [2:0]  st_in_channel,        //       .channel
		output wire [31:0] st_out_data,          // st_out.data
		output wire        st_out_valid,         //       .valid
		input  wire        st_out_ready,         //       .ready
		output wire        st_out_startofpacket, //       .startofpacket
		output wire        st_out_endofpacket,   //       .endofpacket
		output wire [1:0]  st_out_empty,         //       .empty
		output wire [2:0]  st_out_error,         //       .error
		output wire [2:0]  st_out_channel        //       .channel
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (4),
		.BITS_PER_SYMBOL     (8),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (3),
		.ERROR_WIDTH         (3),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dut (
		.clk               (clk_clk),                              //       clk.clk
		.reset             (reset_reset),                          // clk_reset.reset
		.in_data           (st_in_data),                           //        in.data
		.in_valid          (st_in_valid),                          //          .valid
		.in_ready          (st_in_ready),                          //          .ready
		.in_startofpacket  (st_in_startofpacket),                  //          .startofpacket
		.in_endofpacket    (st_in_endofpacket),                    //          .endofpacket
		.in_empty          (st_in_empty),                          //          .empty
		.in_error          (st_in_error),                          //          .error
		.in_channel        (st_in_channel),                        //          .channel
		.out_data          (st_out_data),                          //       out.data
		.out_valid         (st_out_valid),                         //          .valid
		.out_ready         (st_out_ready),                         //          .ready
		.out_startofpacket (st_out_startofpacket),                 //          .startofpacket
		.out_endofpacket   (st_out_endofpacket),                   //          .endofpacket
		.out_empty         (st_out_empty),                         //          .empty
		.out_error         (st_out_error),                         //          .error
		.out_channel       (st_out_channel),                       //          .channel
		.csr_address       (2'b00),                                // (terminated)
		.csr_read          (1'b0),                                 // (terminated)
		.csr_write         (1'b0),                                 // (terminated)
		.csr_readdata      (),                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000), // (terminated)
		.almost_full_data  (),                                     // (terminated)
		.almost_empty_data ()                                      // (terminated)
	);

endmodule
