//----------------------------------------------------------------------------------------------------
// This is the top file of the example test for Avalon Streaming BFM user guide
// The Qsys test bench system and the test program are instantiated.
//----------------------------------------------------------------------------------------------------

module top ();
	st_bfm_qsys_tutorial_tb tb();
	test_program pgm();
endmodule
