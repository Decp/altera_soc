// mityarm_5csx_dev_board.v

// Generated using ACDS version 13.1 162 at 2014.02.17.18:44:51

`timescale 1 ps / 1 ps
module mityarm_5csx_dev_board (
		output wire [14:0] hps_ddr_mem_a,                   // hps_ddr.mem_a
		output wire [2:0]  hps_ddr_mem_ba,                  //        .mem_ba
		output wire        hps_ddr_mem_ck,                  //        .mem_ck
		output wire        hps_ddr_mem_ck_n,                //        .mem_ck_n
		output wire        hps_ddr_mem_cke,                 //        .mem_cke
		output wire        hps_ddr_mem_cs_n,                //        .mem_cs_n
		output wire        hps_ddr_mem_ras_n,               //        .mem_ras_n
		output wire        hps_ddr_mem_cas_n,               //        .mem_cas_n
		output wire        hps_ddr_mem_we_n,                //        .mem_we_n
		output wire        hps_ddr_mem_reset_n,             //        .mem_reset_n
		inout  wire [39:0] hps_ddr_mem_dq,                  //        .mem_dq
		inout  wire [4:0]  hps_ddr_mem_dqs,                 //        .mem_dqs
		inout  wire [4:0]  hps_ddr_mem_dqs_n,               //        .mem_dqs_n
		output wire        hps_ddr_mem_odt,                 //        .mem_odt
		output wire [4:0]  hps_ddr_mem_dm,                  //        .mem_dm
		input  wire        hps_ddr_oct_rzqin,               //        .oct_rzqin
		output wire        hps_io_hps_io_emac1_inst_TX_CLK, //  hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_io_hps_io_emac1_inst_TXD0,   //        .hps_io_emac1_inst_TXD0
		output wire        hps_io_hps_io_emac1_inst_TXD1,   //        .hps_io_emac1_inst_TXD1
		output wire        hps_io_hps_io_emac1_inst_TXD2,   //        .hps_io_emac1_inst_TXD2
		output wire        hps_io_hps_io_emac1_inst_TXD3,   //        .hps_io_emac1_inst_TXD3
		input  wire        hps_io_hps_io_emac1_inst_RXD0,   //        .hps_io_emac1_inst_RXD0
		inout  wire        hps_io_hps_io_emac1_inst_MDIO,   //        .hps_io_emac1_inst_MDIO
		output wire        hps_io_hps_io_emac1_inst_MDC,    //        .hps_io_emac1_inst_MDC
		input  wire        hps_io_hps_io_emac1_inst_RX_CTL, //        .hps_io_emac1_inst_RX_CTL
		output wire        hps_io_hps_io_emac1_inst_TX_CTL, //        .hps_io_emac1_inst_TX_CTL
		input  wire        hps_io_hps_io_emac1_inst_RX_CLK, //        .hps_io_emac1_inst_RX_CLK
		input  wire        hps_io_hps_io_emac1_inst_RXD1,   //        .hps_io_emac1_inst_RXD1
		input  wire        hps_io_hps_io_emac1_inst_RXD2,   //        .hps_io_emac1_inst_RXD2
		input  wire        hps_io_hps_io_emac1_inst_RXD3,   //        .hps_io_emac1_inst_RXD3
		output wire        hps_io_hps_io_qspi_inst_SS1,     //        .hps_io_qspi_inst_SS1
		inout  wire        hps_io_hps_io_qspi_inst_IO0,     //        .hps_io_qspi_inst_IO0
		inout  wire        hps_io_hps_io_qspi_inst_IO1,     //        .hps_io_qspi_inst_IO1
		inout  wire        hps_io_hps_io_qspi_inst_IO2,     //        .hps_io_qspi_inst_IO2
		inout  wire        hps_io_hps_io_qspi_inst_IO3,     //        .hps_io_qspi_inst_IO3
		output wire        hps_io_hps_io_qspi_inst_SS0,     //        .hps_io_qspi_inst_SS0
		output wire        hps_io_hps_io_qspi_inst_CLK,     //        .hps_io_qspi_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_CMD,     //        .hps_io_sdio_inst_CMD
		inout  wire        hps_io_hps_io_sdio_inst_D0,      //        .hps_io_sdio_inst_D0
		inout  wire        hps_io_hps_io_sdio_inst_D1,      //        .hps_io_sdio_inst_D1
		output wire        hps_io_hps_io_sdio_inst_CLK,     //        .hps_io_sdio_inst_CLK
		inout  wire        hps_io_hps_io_sdio_inst_D2,      //        .hps_io_sdio_inst_D2
		inout  wire        hps_io_hps_io_sdio_inst_D3,      //        .hps_io_sdio_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D0,      //        .hps_io_usb1_inst_D0
		inout  wire        hps_io_hps_io_usb1_inst_D1,      //        .hps_io_usb1_inst_D1
		inout  wire        hps_io_hps_io_usb1_inst_D2,      //        .hps_io_usb1_inst_D2
		inout  wire        hps_io_hps_io_usb1_inst_D3,      //        .hps_io_usb1_inst_D3
		inout  wire        hps_io_hps_io_usb1_inst_D4,      //        .hps_io_usb1_inst_D4
		inout  wire        hps_io_hps_io_usb1_inst_D5,      //        .hps_io_usb1_inst_D5
		inout  wire        hps_io_hps_io_usb1_inst_D6,      //        .hps_io_usb1_inst_D6
		inout  wire        hps_io_hps_io_usb1_inst_D7,      //        .hps_io_usb1_inst_D7
		input  wire        hps_io_hps_io_usb1_inst_CLK,     //        .hps_io_usb1_inst_CLK
		output wire        hps_io_hps_io_usb1_inst_STP,     //        .hps_io_usb1_inst_STP
		input  wire        hps_io_hps_io_usb1_inst_DIR,     //        .hps_io_usb1_inst_DIR
		input  wire        hps_io_hps_io_usb1_inst_NXT,     //        .hps_io_usb1_inst_NXT
		input  wire        hps_io_hps_io_uart0_inst_RX,     //        .hps_io_uart0_inst_RX
		output wire        hps_io_hps_io_uart0_inst_TX,     //        .hps_io_uart0_inst_TX
		inout  wire        hps_io_hps_io_i2c0_inst_SDA,     //        .hps_io_i2c0_inst_SDA
		inout  wire        hps_io_hps_io_i2c0_inst_SCL,     //        .hps_io_i2c0_inst_SCL
		inout  wire        hps_io_hps_io_i2c1_inst_SDA,     //        .hps_io_i2c1_inst_SDA
		inout  wire        hps_io_hps_io_i2c1_inst_SCL,     //        .hps_io_i2c1_inst_SCL
		input  wire        hps_io_hps_io_can0_inst_RX,      //        .hps_io_can0_inst_RX
		output wire        hps_io_hps_io_can0_inst_TX,      //        .hps_io_can0_inst_TX
		input  wire        hps_io_hps_io_can1_inst_RX,      //        .hps_io_can1_inst_RX
		output wire        hps_io_hps_io_can1_inst_TX,      //        .hps_io_can1_inst_TX
		inout  wire        hps_io_hps_io_gpio_inst_GPIO00,  //        .hps_io_gpio_inst_GPIO00
		inout  wire        hps_io_hps_io_gpio_inst_GPIO09,  //        .hps_io_gpio_inst_GPIO09
		inout  wire        hps_io_hps_io_gpio_inst_GPIO28,  //        .hps_io_gpio_inst_GPIO28
		inout  wire        hps_io_hps_io_gpio_inst_GPIO37,  //        .hps_io_gpio_inst_GPIO37
		inout  wire        hps_io_hps_io_gpio_inst_GPIO40,  //        .hps_io_gpio_inst_GPIO40
		inout  wire        hps_io_hps_io_gpio_inst_GPIO41,  //        .hps_io_gpio_inst_GPIO41
		inout  wire        hps_io_hps_io_gpio_inst_GPIO48,  //        .hps_io_gpio_inst_GPIO48
		inout  wire        hps_io_hps_io_gpio_inst_GPIO49,  //        .hps_io_gpio_inst_GPIO49
		inout  wire        hps_io_hps_io_gpio_inst_GPIO50   //        .hps_io_gpio_inst_GPIO50
	);

	wire          hps_0_h2f_user0_clock_clk;                                                 // hps_0:h2f_user0_clk -> [dma_write_master_0:clk, hps_0:f2h_sdram0_clk, hps_0:h2f_lw_axi_clk, mm_interconnect_0:hps_0_h2f_user0_clock_clk, mm_interconnect_1:hps_0_h2f_user0_clock_clk, modular_sgdma_dispatcher_0:clk, rst_controller:clk, sysid_qsys:clock]
	wire          modular_sgdma_dispatcher_0_write_command_source_valid;                     // modular_sgdma_dispatcher_0:src_write_master_valid -> dma_write_master_0:snk_command_valid
	wire  [255:0] modular_sgdma_dispatcher_0_write_command_source_data;                      // modular_sgdma_dispatcher_0:src_write_master_data -> dma_write_master_0:snk_command_data
	wire          modular_sgdma_dispatcher_0_write_command_source_ready;                     // dma_write_master_0:snk_command_ready -> modular_sgdma_dispatcher_0:src_write_master_ready
	wire          dma_write_master_0_response_source_valid;                                  // dma_write_master_0:src_response_valid -> modular_sgdma_dispatcher_0:snk_write_master_valid
	wire  [255:0] dma_write_master_0_response_source_data;                                   // dma_write_master_0:src_response_data -> modular_sgdma_dispatcher_0:snk_write_master_data
	wire          dma_write_master_0_response_source_ready;                                  // modular_sgdma_dispatcher_0:snk_write_master_ready -> dma_write_master_0:src_response_ready
	wire    [0:0] mm_interconnect_0_sysid_qsys_control_slave_address;                        // mm_interconnect_0:sysid_qsys_control_slave_address -> sysid_qsys:address
	wire   [31:0] mm_interconnect_0_sysid_qsys_control_slave_readdata;                       // sysid_qsys:readdata -> mm_interconnect_0:sysid_qsys_control_slave_readdata
	wire          mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_waitrequest; // modular_sgdma_dispatcher_0:descriptor_waitrequest -> mm_interconnect_0:modular_sgdma_dispatcher_0_Descriptor_Slave_waitrequest
	wire  [127:0] mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_writedata;   // mm_interconnect_0:modular_sgdma_dispatcher_0_Descriptor_Slave_writedata -> modular_sgdma_dispatcher_0:descriptor_writedata
	wire          mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_write;       // mm_interconnect_0:modular_sgdma_dispatcher_0_Descriptor_Slave_write -> modular_sgdma_dispatcher_0:descriptor_write
	wire   [15:0] mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_byteenable;  // mm_interconnect_0:modular_sgdma_dispatcher_0_Descriptor_Slave_byteenable -> modular_sgdma_dispatcher_0:descriptor_byteenable
	wire   [31:0] mm_interconnect_0_modular_sgdma_dispatcher_0_csr_writedata;                // mm_interconnect_0:modular_sgdma_dispatcher_0_CSR_writedata -> modular_sgdma_dispatcher_0:csr_writedata
	wire    [2:0] mm_interconnect_0_modular_sgdma_dispatcher_0_csr_address;                  // mm_interconnect_0:modular_sgdma_dispatcher_0_CSR_address -> modular_sgdma_dispatcher_0:csr_address
	wire          mm_interconnect_0_modular_sgdma_dispatcher_0_csr_write;                    // mm_interconnect_0:modular_sgdma_dispatcher_0_CSR_write -> modular_sgdma_dispatcher_0:csr_write
	wire          mm_interconnect_0_modular_sgdma_dispatcher_0_csr_read;                     // mm_interconnect_0:modular_sgdma_dispatcher_0_CSR_read -> modular_sgdma_dispatcher_0:csr_read
	wire   [31:0] mm_interconnect_0_modular_sgdma_dispatcher_0_csr_readdata;                 // modular_sgdma_dispatcher_0:csr_readdata -> mm_interconnect_0:modular_sgdma_dispatcher_0_CSR_readdata
	wire    [3:0] mm_interconnect_0_modular_sgdma_dispatcher_0_csr_byteenable;               // mm_interconnect_0:modular_sgdma_dispatcher_0_CSR_byteenable -> modular_sgdma_dispatcher_0:csr_byteenable
	wire          hps_0_h2f_lw_axi_master_awvalid;                                           // hps_0:h2f_lw_AWVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                            // hps_0:h2f_lw_ARSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arsize
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                            // hps_0:h2f_lw_ARLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlock
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                           // hps_0:h2f_lw_AWCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awcache
	wire          hps_0_h2f_lw_axi_master_arready;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_arready -> hps_0:h2f_lw_ARREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                              // hps_0:h2f_lw_ARID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arid
	wire          hps_0_h2f_lw_axi_master_rready;                                            // hps_0:h2f_lw_RREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_rready
	wire          hps_0_h2f_lw_axi_master_bready;                                            // hps_0:h2f_lw_BREADY -> mm_interconnect_0:hps_0_h2f_lw_axi_master_bready
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                            // hps_0:h2f_lw_AWSIZE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awsize
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                            // hps_0:h2f_lw_AWPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awprot
	wire          hps_0_h2f_lw_axi_master_arvalid;                                           // hps_0:h2f_lw_ARVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                            // hps_0:h2f_lw_ARPROT -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arprot
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_bid -> hps_0:h2f_lw_BID
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                             // hps_0:h2f_lw_ARLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arlen
	wire          hps_0_h2f_lw_axi_master_awready;                                           // mm_interconnect_0:hps_0_h2f_lw_axi_master_awready -> hps_0:h2f_lw_AWREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                              // hps_0:h2f_lw_AWID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awid
	wire          hps_0_h2f_lw_axi_master_bvalid;                                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_bvalid -> hps_0:h2f_lw_BVALID
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                               // hps_0:h2f_lw_WID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wid
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                            // hps_0:h2f_lw_AWLOCK -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                           // hps_0:h2f_lw_AWBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awburst
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_bresp -> hps_0:h2f_lw_BRESP
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                             // hps_0:h2f_lw_WSTRB -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wstrb
	wire          hps_0_h2f_lw_axi_master_rvalid;                                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                             // hps_0:h2f_lw_WDATA -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wdata
	wire          hps_0_h2f_lw_axi_master_wready;                                            // mm_interconnect_0:hps_0_h2f_lw_axi_master_wready -> hps_0:h2f_lw_WREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                           // hps_0:h2f_lw_ARBURST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arburst
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rdata -> hps_0:h2f_lw_RDATA
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                            // hps_0:h2f_lw_ARADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_araddr
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                           // hps_0:h2f_lw_ARCACHE -> mm_interconnect_0:hps_0_h2f_lw_axi_master_arcache
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                             // hps_0:h2f_lw_AWLEN -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awlen
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                            // hps_0:h2f_lw_AWADDR -> mm_interconnect_0:hps_0_h2f_lw_axi_master_awaddr
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                               // mm_interconnect_0:hps_0_h2f_lw_axi_master_rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_wvalid;                                            // hps_0:h2f_lw_WVALID -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wvalid
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rresp -> hps_0:h2f_lw_RRESP
	wire          hps_0_h2f_lw_axi_master_wlast;                                             // hps_0:h2f_lw_WLAST -> mm_interconnect_0:hps_0_h2f_lw_axi_master_wlast
	wire          hps_0_h2f_lw_axi_master_rlast;                                             // mm_interconnect_0:hps_0_h2f_lw_axi_master_rlast -> hps_0:h2f_lw_RLAST
	wire    [5:0] dma_write_master_0_data_write_master_burstcount;                           // dma_write_master_0:master_burstcount -> mm_interconnect_1:dma_write_master_0_Data_Write_Master_burstcount
	wire          dma_write_master_0_data_write_master_waitrequest;                          // mm_interconnect_1:dma_write_master_0_Data_Write_Master_waitrequest -> dma_write_master_0:master_waitrequest
	wire   [63:0] dma_write_master_0_data_write_master_writedata;                            // dma_write_master_0:master_writedata -> mm_interconnect_1:dma_write_master_0_Data_Write_Master_writedata
	wire   [31:0] dma_write_master_0_data_write_master_address;                              // dma_write_master_0:master_address -> mm_interconnect_1:dma_write_master_0_Data_Write_Master_address
	wire          dma_write_master_0_data_write_master_write;                                // dma_write_master_0:master_write -> mm_interconnect_1:dma_write_master_0_Data_Write_Master_write
	wire    [7:0] dma_write_master_0_data_write_master_byteenable;                           // dma_write_master_0:master_byteenable -> mm_interconnect_1:dma_write_master_0_Data_Write_Master_byteenable
	wire          mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest;                       // hps_0:f2h_sdram0_WAITREQUEST -> mm_interconnect_1:hps_0_f2h_sdram0_data_waitrequest
	wire    [7:0] mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount;                        // mm_interconnect_1:hps_0_f2h_sdram0_data_burstcount -> hps_0:f2h_sdram0_BURSTCOUNT
	wire   [63:0] mm_interconnect_1_hps_0_f2h_sdram0_data_writedata;                         // mm_interconnect_1:hps_0_f2h_sdram0_data_writedata -> hps_0:f2h_sdram0_WRITEDATA
	wire   [28:0] mm_interconnect_1_hps_0_f2h_sdram0_data_address;                           // mm_interconnect_1:hps_0_f2h_sdram0_data_address -> hps_0:f2h_sdram0_ADDRESS
	wire          mm_interconnect_1_hps_0_f2h_sdram0_data_write;                             // mm_interconnect_1:hps_0_f2h_sdram0_data_write -> hps_0:f2h_sdram0_WRITE
	wire    [7:0] mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable;                        // mm_interconnect_1:hps_0_f2h_sdram0_data_byteenable -> hps_0:f2h_sdram0_BYTEENABLE
	wire   [31:0] hps_0_f2h_irq0_irq;                                                        // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                        // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          rst_controller_reset_out_reset;                                            // rst_controller:reset_out -> [dma_write_master_0:reset, mm_interconnect_0:sysid_qsys_reset_reset_bridge_in_reset_reset, mm_interconnect_1:dma_write_master_0_Clock_reset_reset_bridge_in_reset_reset, modular_sgdma_dispatcher_0:reset, sysid_qsys:reset_n]
	wire          hps_0_h2f_reset_reset;                                                     // hps_0:h2f_rst_n -> rst_controller:reset_in0

	mityarm_5csx_dev_board_hps_0 #(
		.F2S_Width (0),
		.S2F_Width (0)
	) hps_0 (
		.h2f_user0_clk            (hps_0_h2f_user0_clock_clk),                           //   h2f_user0_clock.clk
		.mem_a                    (hps_ddr_mem_a),                                       //            memory.mem_a
		.mem_ba                   (hps_ddr_mem_ba),                                      //                  .mem_ba
		.mem_ck                   (hps_ddr_mem_ck),                                      //                  .mem_ck
		.mem_ck_n                 (hps_ddr_mem_ck_n),                                    //                  .mem_ck_n
		.mem_cke                  (hps_ddr_mem_cke),                                     //                  .mem_cke
		.mem_cs_n                 (hps_ddr_mem_cs_n),                                    //                  .mem_cs_n
		.mem_ras_n                (hps_ddr_mem_ras_n),                                   //                  .mem_ras_n
		.mem_cas_n                (hps_ddr_mem_cas_n),                                   //                  .mem_cas_n
		.mem_we_n                 (hps_ddr_mem_we_n),                                    //                  .mem_we_n
		.mem_reset_n              (hps_ddr_mem_reset_n),                                 //                  .mem_reset_n
		.mem_dq                   (hps_ddr_mem_dq),                                      //                  .mem_dq
		.mem_dqs                  (hps_ddr_mem_dqs),                                     //                  .mem_dqs
		.mem_dqs_n                (hps_ddr_mem_dqs_n),                                   //                  .mem_dqs_n
		.mem_odt                  (hps_ddr_mem_odt),                                     //                  .mem_odt
		.mem_dm                   (hps_ddr_mem_dm),                                      //                  .mem_dm
		.oct_rzqin                (hps_ddr_oct_rzqin),                                   //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_io_hps_io_emac1_inst_TX_CLK),                     //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_io_hps_io_emac1_inst_TXD0),                       //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_io_hps_io_emac1_inst_TXD1),                       //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_io_hps_io_emac1_inst_TXD2),                       //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_io_hps_io_emac1_inst_TXD3),                       //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_io_hps_io_emac1_inst_RXD0),                       //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_io_hps_io_emac1_inst_MDIO),                       //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_io_hps_io_emac1_inst_MDC),                        //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_io_hps_io_emac1_inst_RX_CTL),                     //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_io_hps_io_emac1_inst_TX_CTL),                     //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_io_hps_io_emac1_inst_RX_CLK),                     //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_io_hps_io_emac1_inst_RXD1),                       //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_io_hps_io_emac1_inst_RXD2),                       //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_io_hps_io_emac1_inst_RXD3),                       //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_SS1     (hps_io_hps_io_qspi_inst_SS1),                         //                  .hps_io_qspi_inst_SS1
		.hps_io_qspi_inst_IO0     (hps_io_hps_io_qspi_inst_IO0),                         //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_io_hps_io_qspi_inst_IO1),                         //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_io_hps_io_qspi_inst_IO2),                         //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_io_hps_io_qspi_inst_IO3),                         //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_io_hps_io_qspi_inst_SS0),                         //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_io_hps_io_qspi_inst_CLK),                         //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_io_hps_io_sdio_inst_CMD),                         //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_io_hps_io_sdio_inst_D0),                          //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_io_hps_io_sdio_inst_D1),                          //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_io_hps_io_sdio_inst_CLK),                         //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_io_hps_io_sdio_inst_D2),                          //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_io_hps_io_sdio_inst_D3),                          //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_io_hps_io_usb1_inst_D0),                          //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_io_hps_io_usb1_inst_D1),                          //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_io_hps_io_usb1_inst_D2),                          //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_io_hps_io_usb1_inst_D3),                          //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_io_hps_io_usb1_inst_D4),                          //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_io_hps_io_usb1_inst_D5),                          //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_io_hps_io_usb1_inst_D6),                          //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_io_hps_io_usb1_inst_D7),                          //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_io_hps_io_usb1_inst_CLK),                         //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_io_hps_io_usb1_inst_STP),                         //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_io_hps_io_usb1_inst_DIR),                         //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_io_hps_io_usb1_inst_NXT),                         //                  .hps_io_usb1_inst_NXT
		.hps_io_uart0_inst_RX     (hps_io_hps_io_uart0_inst_RX),                         //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_io_hps_io_uart0_inst_TX),                         //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_io_hps_io_i2c0_inst_SDA),                         //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_io_hps_io_i2c0_inst_SCL),                         //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_io_hps_io_i2c1_inst_SDA),                         //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_io_hps_io_i2c1_inst_SCL),                         //                  .hps_io_i2c1_inst_SCL
		.hps_io_can0_inst_RX      (hps_io_hps_io_can0_inst_RX),                          //                  .hps_io_can0_inst_RX
		.hps_io_can0_inst_TX      (hps_io_hps_io_can0_inst_TX),                          //                  .hps_io_can0_inst_TX
		.hps_io_can1_inst_RX      (hps_io_hps_io_can1_inst_RX),                          //                  .hps_io_can1_inst_RX
		.hps_io_can1_inst_TX      (hps_io_hps_io_can1_inst_TX),                          //                  .hps_io_can1_inst_TX
		.hps_io_gpio_inst_GPIO00  (hps_io_hps_io_gpio_inst_GPIO00),                      //                  .hps_io_gpio_inst_GPIO00
		.hps_io_gpio_inst_GPIO09  (hps_io_hps_io_gpio_inst_GPIO09),                      //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO28  (hps_io_hps_io_gpio_inst_GPIO28),                      //                  .hps_io_gpio_inst_GPIO28
		.hps_io_gpio_inst_GPIO37  (hps_io_hps_io_gpio_inst_GPIO37),                      //                  .hps_io_gpio_inst_GPIO37
		.hps_io_gpio_inst_GPIO40  (hps_io_hps_io_gpio_inst_GPIO40),                      //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_io_hps_io_gpio_inst_GPIO41),                      //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_io_hps_io_gpio_inst_GPIO48),                      //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO49  (hps_io_hps_io_gpio_inst_GPIO49),                      //                  .hps_io_gpio_inst_GPIO49
		.hps_io_gpio_inst_GPIO50  (hps_io_hps_io_gpio_inst_GPIO50),                      //                  .hps_io_gpio_inst_GPIO50
		.h2f_rst_n                (hps_0_h2f_reset_reset),                               //         h2f_reset.reset_n
		.f2h_sdram0_clk           (hps_0_h2f_user0_clock_clk),                           //  f2h_sdram0_clock.clk
		.f2h_sdram0_ADDRESS       (mm_interconnect_1_hps_0_f2h_sdram0_data_address),     //   f2h_sdram0_data.address
		.f2h_sdram0_BURSTCOUNT    (mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount),  //                  .burstcount
		.f2h_sdram0_WAITREQUEST   (mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest), //                  .waitrequest
		.f2h_sdram0_WRITEDATA     (mm_interconnect_1_hps_0_f2h_sdram0_data_writedata),   //                  .writedata
		.f2h_sdram0_BYTEENABLE    (mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable),  //                  .byteenable
		.f2h_sdram0_WRITE         (mm_interconnect_1_hps_0_f2h_sdram0_data_write),       //                  .write
		.h2f_lw_axi_clk           (hps_0_h2f_user0_clock_clk),                           //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                        // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                      //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                       //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                      //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                     //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                      //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                     //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                      //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                     //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                     //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                         //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                       //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                       //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                       //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                      //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                      //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                         //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                       //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                      //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                      //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                        //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                      //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                       //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                      //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                     //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                      //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                     //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                      //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                     //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                     //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                         //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                       //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                       //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                       //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                      //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                      //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                                  //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                                   //          f2h_irq1.irq
	);

	mityarm_5csx_dev_board_sysid_qsys sysid_qsys (
		.clock    (hps_0_h2f_user0_clock_clk),                           //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                     //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_qsys_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_qsys_control_slave_address)   //              .address
	);

	dispatcher #(
		.MODE                        (2),
		.RESPONSE_PORT               (2),
		.DESCRIPTOR_FIFO_DEPTH       (8),
		.ENHANCED_FEATURES           (0),
		.DESCRIPTOR_WIDTH            (128),
		.DESCRIPTOR_BYTEENABLE_WIDTH (16),
		.CSR_ADDRESS_WIDTH           (3)
	) modular_sgdma_dispatcher_0 (
		.clk                     (hps_0_h2f_user0_clock_clk),                                                                                                                                                                                                                                             //                clock.clk
		.reset                   (rst_controller_reset_out_reset),                                                                                                                                                                                                                                        //          clock_reset.reset
		.csr_writedata           (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_writedata),                                                                                                                                                                                                            //                  CSR.writedata
		.csr_write               (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_write),                                                                                                                                                                                                                //                     .write
		.csr_byteenable          (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_byteenable),                                                                                                                                                                                                           //                     .byteenable
		.csr_readdata            (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_readdata),                                                                                                                                                                                                             //                     .readdata
		.csr_read                (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_read),                                                                                                                                                                                                                 //                     .read
		.csr_address             (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_address),                                                                                                                                                                                                              //                     .address
		.descriptor_write        (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_write),                                                                                                                                                                                                   //     Descriptor_Slave.write
		.descriptor_waitrequest  (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_waitrequest),                                                                                                                                                                                             //                     .waitrequest
		.descriptor_writedata    (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_writedata),                                                                                                                                                                                               //                     .writedata
		.descriptor_byteenable   (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_byteenable),                                                                                                                                                                                              //                     .byteenable
		.src_write_master_data   (modular_sgdma_dispatcher_0_write_command_source_data),                                                                                                                                                                                                                  // Write_Command_Source.data
		.src_write_master_valid  (modular_sgdma_dispatcher_0_write_command_source_valid),                                                                                                                                                                                                                 //                     .valid
		.src_write_master_ready  (modular_sgdma_dispatcher_0_write_command_source_ready),                                                                                                                                                                                                                 //                     .ready
		.snk_write_master_data   (dma_write_master_0_response_source_data),                                                                                                                                                                                                                               //  Write_Response_Sink.data
		.snk_write_master_valid  (dma_write_master_0_response_source_valid),                                                                                                                                                                                                                              //                     .valid
		.snk_write_master_ready  (dma_write_master_0_response_source_ready),                                                                                                                                                                                                                              //                     .ready
		.csr_irq                 (),                                                                                                                                                                                                                                                                      //              csr_irq.irq
		.src_response_data       (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_response_valid      (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_response_ready      (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.mm_response_waitrequest (),                                                                                                                                                                                                                                                                      //          (terminated)
		.mm_response_byteenable  (4'b0000),                                                                                                                                                                                                                                                               //          (terminated)
		.mm_response_address     (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.mm_response_readdata    (),                                                                                                                                                                                                                                                                      //          (terminated)
		.mm_response_read        (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.src_read_master_data    (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_read_master_valid   (),                                                                                                                                                                                                                                                                      //          (terminated)
		.src_read_master_ready   (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.snk_read_master_data    (256'b0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000), //          (terminated)
		.snk_read_master_valid   (1'b0),                                                                                                                                                                                                                                                                  //          (terminated)
		.snk_read_master_ready   ()                                                                                                                                                                                                                                                                       //          (terminated)
	);

	write_master #(
		.DATA_WIDTH                     (64),
		.LENGTH_WIDTH                   (32),
		.FIFO_DEPTH                     (128),
		.STRIDE_ENABLE                  (0),
		.BURST_ENABLE                   (1),
		.PACKET_ENABLE                  (1),
		.ERROR_ENABLE                   (0),
		.ERROR_WIDTH                    (8),
		.BYTE_ENABLE_WIDTH              (8),
		.BYTE_ENABLE_WIDTH_LOG2         (3),
		.ADDRESS_WIDTH                  (32),
		.FIFO_DEPTH_LOG2                (7),
		.SYMBOL_WIDTH                   (8),
		.NUMBER_OF_SYMBOLS              (8),
		.NUMBER_OF_SYMBOLS_LOG2         (3),
		.MAX_BURST_COUNT_WIDTH          (6),
		.UNALIGNED_ACCESSES_ENABLE      (0),
		.ONLY_FULL_ACCESS_ENABLE        (0),
		.BURST_WRAPPING_SUPPORT         (0),
		.PROGRAMMABLE_BURST_ENABLE      (0),
		.MAX_BURST_COUNT                (32),
		.FIFO_SPEED_OPTIMIZATION        (1),
		.STRIDE_WIDTH                   (1),
		.ACTUAL_BYTES_TRANSFERRED_WIDTH (32)
	) dma_write_master_0 (
		.clk                (hps_0_h2f_user0_clock_clk),                             //             Clock.clk
		.reset              (rst_controller_reset_out_reset),                        //       Clock_reset.reset
		.master_address     (dma_write_master_0_data_write_master_address),          // Data_Write_Master.address
		.master_write       (dma_write_master_0_data_write_master_write),            //                  .write
		.master_byteenable  (dma_write_master_0_data_write_master_byteenable),       //                  .byteenable
		.master_writedata   (dma_write_master_0_data_write_master_writedata),        //                  .writedata
		.master_waitrequest (dma_write_master_0_data_write_master_waitrequest),      //                  .waitrequest
		.master_burstcount  (dma_write_master_0_data_write_master_burstcount),       //                  .burstcount
		.snk_data           (),                                                      //         Data_Sink.data
		.snk_valid          (),                                                      //                  .valid
		.snk_ready          (),                                                      //                  .ready
		.snk_sop            (),                                                      //                  .startofpacket
		.snk_eop            (),                                                      //                  .endofpacket
		.snk_empty          (),                                                      //                  .empty
		.snk_command_data   (modular_sgdma_dispatcher_0_write_command_source_data),  //      Command_Sink.data
		.snk_command_valid  (modular_sgdma_dispatcher_0_write_command_source_valid), //                  .valid
		.snk_command_ready  (modular_sgdma_dispatcher_0_write_command_source_ready), //                  .ready
		.src_response_data  (dma_write_master_0_response_source_data),               //   Response_Source.data
		.src_response_valid (dma_write_master_0_response_source_valid),              //                  .valid
		.src_response_ready (dma_write_master_0_response_source_ready),              //                  .ready
		.snk_error          (8'b00000000)                                            //       (terminated)
	);

	mityarm_5csx_dev_board_mm_interconnect_0 mm_interconnect_0 (
		.hps_0_h2f_lw_axi_master_awid                            (hps_0_h2f_lw_axi_master_awid),                                              //                     hps_0_h2f_lw_axi_master.awid
		.hps_0_h2f_lw_axi_master_awaddr                          (hps_0_h2f_lw_axi_master_awaddr),                                            //                                            .awaddr
		.hps_0_h2f_lw_axi_master_awlen                           (hps_0_h2f_lw_axi_master_awlen),                                             //                                            .awlen
		.hps_0_h2f_lw_axi_master_awsize                          (hps_0_h2f_lw_axi_master_awsize),                                            //                                            .awsize
		.hps_0_h2f_lw_axi_master_awburst                         (hps_0_h2f_lw_axi_master_awburst),                                           //                                            .awburst
		.hps_0_h2f_lw_axi_master_awlock                          (hps_0_h2f_lw_axi_master_awlock),                                            //                                            .awlock
		.hps_0_h2f_lw_axi_master_awcache                         (hps_0_h2f_lw_axi_master_awcache),                                           //                                            .awcache
		.hps_0_h2f_lw_axi_master_awprot                          (hps_0_h2f_lw_axi_master_awprot),                                            //                                            .awprot
		.hps_0_h2f_lw_axi_master_awvalid                         (hps_0_h2f_lw_axi_master_awvalid),                                           //                                            .awvalid
		.hps_0_h2f_lw_axi_master_awready                         (hps_0_h2f_lw_axi_master_awready),                                           //                                            .awready
		.hps_0_h2f_lw_axi_master_wid                             (hps_0_h2f_lw_axi_master_wid),                                               //                                            .wid
		.hps_0_h2f_lw_axi_master_wdata                           (hps_0_h2f_lw_axi_master_wdata),                                             //                                            .wdata
		.hps_0_h2f_lw_axi_master_wstrb                           (hps_0_h2f_lw_axi_master_wstrb),                                             //                                            .wstrb
		.hps_0_h2f_lw_axi_master_wlast                           (hps_0_h2f_lw_axi_master_wlast),                                             //                                            .wlast
		.hps_0_h2f_lw_axi_master_wvalid                          (hps_0_h2f_lw_axi_master_wvalid),                                            //                                            .wvalid
		.hps_0_h2f_lw_axi_master_wready                          (hps_0_h2f_lw_axi_master_wready),                                            //                                            .wready
		.hps_0_h2f_lw_axi_master_bid                             (hps_0_h2f_lw_axi_master_bid),                                               //                                            .bid
		.hps_0_h2f_lw_axi_master_bresp                           (hps_0_h2f_lw_axi_master_bresp),                                             //                                            .bresp
		.hps_0_h2f_lw_axi_master_bvalid                          (hps_0_h2f_lw_axi_master_bvalid),                                            //                                            .bvalid
		.hps_0_h2f_lw_axi_master_bready                          (hps_0_h2f_lw_axi_master_bready),                                            //                                            .bready
		.hps_0_h2f_lw_axi_master_arid                            (hps_0_h2f_lw_axi_master_arid),                                              //                                            .arid
		.hps_0_h2f_lw_axi_master_araddr                          (hps_0_h2f_lw_axi_master_araddr),                                            //                                            .araddr
		.hps_0_h2f_lw_axi_master_arlen                           (hps_0_h2f_lw_axi_master_arlen),                                             //                                            .arlen
		.hps_0_h2f_lw_axi_master_arsize                          (hps_0_h2f_lw_axi_master_arsize),                                            //                                            .arsize
		.hps_0_h2f_lw_axi_master_arburst                         (hps_0_h2f_lw_axi_master_arburst),                                           //                                            .arburst
		.hps_0_h2f_lw_axi_master_arlock                          (hps_0_h2f_lw_axi_master_arlock),                                            //                                            .arlock
		.hps_0_h2f_lw_axi_master_arcache                         (hps_0_h2f_lw_axi_master_arcache),                                           //                                            .arcache
		.hps_0_h2f_lw_axi_master_arprot                          (hps_0_h2f_lw_axi_master_arprot),                                            //                                            .arprot
		.hps_0_h2f_lw_axi_master_arvalid                         (hps_0_h2f_lw_axi_master_arvalid),                                           //                                            .arvalid
		.hps_0_h2f_lw_axi_master_arready                         (hps_0_h2f_lw_axi_master_arready),                                           //                                            .arready
		.hps_0_h2f_lw_axi_master_rid                             (hps_0_h2f_lw_axi_master_rid),                                               //                                            .rid
		.hps_0_h2f_lw_axi_master_rdata                           (hps_0_h2f_lw_axi_master_rdata),                                             //                                            .rdata
		.hps_0_h2f_lw_axi_master_rresp                           (hps_0_h2f_lw_axi_master_rresp),                                             //                                            .rresp
		.hps_0_h2f_lw_axi_master_rlast                           (hps_0_h2f_lw_axi_master_rlast),                                             //                                            .rlast
		.hps_0_h2f_lw_axi_master_rvalid                          (hps_0_h2f_lw_axi_master_rvalid),                                            //                                            .rvalid
		.hps_0_h2f_lw_axi_master_rready                          (hps_0_h2f_lw_axi_master_rready),                                            //                                            .rready
		.hps_0_h2f_user0_clock_clk                               (hps_0_h2f_user0_clock_clk),                                                 //                       hps_0_h2f_user0_clock.clk
		.sysid_qsys_reset_reset_bridge_in_reset_reset            (rst_controller_reset_out_reset),                                            //      sysid_qsys_reset_reset_bridge_in_reset.reset
		.modular_sgdma_dispatcher_0_CSR_address                  (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_address),                  //              modular_sgdma_dispatcher_0_CSR.address
		.modular_sgdma_dispatcher_0_CSR_write                    (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_write),                    //                                            .write
		.modular_sgdma_dispatcher_0_CSR_read                     (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_read),                     //                                            .read
		.modular_sgdma_dispatcher_0_CSR_readdata                 (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_readdata),                 //                                            .readdata
		.modular_sgdma_dispatcher_0_CSR_writedata                (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_writedata),                //                                            .writedata
		.modular_sgdma_dispatcher_0_CSR_byteenable               (mm_interconnect_0_modular_sgdma_dispatcher_0_csr_byteenable),               //                                            .byteenable
		.modular_sgdma_dispatcher_0_Descriptor_Slave_write       (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_write),       // modular_sgdma_dispatcher_0_Descriptor_Slave.write
		.modular_sgdma_dispatcher_0_Descriptor_Slave_writedata   (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_writedata),   //                                            .writedata
		.modular_sgdma_dispatcher_0_Descriptor_Slave_byteenable  (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_byteenable),  //                                            .byteenable
		.modular_sgdma_dispatcher_0_Descriptor_Slave_waitrequest (mm_interconnect_0_modular_sgdma_dispatcher_0_descriptor_slave_waitrequest), //                                            .waitrequest
		.sysid_qsys_control_slave_address                        (mm_interconnect_0_sysid_qsys_control_slave_address),                        //                    sysid_qsys_control_slave.address
		.sysid_qsys_control_slave_readdata                       (mm_interconnect_0_sysid_qsys_control_slave_readdata)                        //                                            .readdata
	);

	mityarm_5csx_dev_board_mm_interconnect_1 mm_interconnect_1 (
		.hps_0_h2f_user0_clock_clk                                  (hps_0_h2f_user0_clock_clk),                           //                                hps_0_h2f_user0_clock.clk
		.dma_write_master_0_Clock_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                      // dma_write_master_0_Clock_reset_reset_bridge_in_reset.reset
		.dma_write_master_0_Data_Write_Master_address               (dma_write_master_0_data_write_master_address),        //                 dma_write_master_0_Data_Write_Master.address
		.dma_write_master_0_Data_Write_Master_waitrequest           (dma_write_master_0_data_write_master_waitrequest),    //                                                     .waitrequest
		.dma_write_master_0_Data_Write_Master_burstcount            (dma_write_master_0_data_write_master_burstcount),     //                                                     .burstcount
		.dma_write_master_0_Data_Write_Master_byteenable            (dma_write_master_0_data_write_master_byteenable),     //                                                     .byteenable
		.dma_write_master_0_Data_Write_Master_write                 (dma_write_master_0_data_write_master_write),          //                                                     .write
		.dma_write_master_0_Data_Write_Master_writedata             (dma_write_master_0_data_write_master_writedata),      //                                                     .writedata
		.hps_0_f2h_sdram0_data_address                              (mm_interconnect_1_hps_0_f2h_sdram0_data_address),     //                                hps_0_f2h_sdram0_data.address
		.hps_0_f2h_sdram0_data_write                                (mm_interconnect_1_hps_0_f2h_sdram0_data_write),       //                                                     .write
		.hps_0_f2h_sdram0_data_writedata                            (mm_interconnect_1_hps_0_f2h_sdram0_data_writedata),   //                                                     .writedata
		.hps_0_f2h_sdram0_data_burstcount                           (mm_interconnect_1_hps_0_f2h_sdram0_data_burstcount),  //                                                     .burstcount
		.hps_0_f2h_sdram0_data_byteenable                           (mm_interconnect_1_hps_0_f2h_sdram0_data_byteenable),  //                                                     .byteenable
		.hps_0_f2h_sdram0_data_waitrequest                          (mm_interconnect_1_hps_0_f2h_sdram0_data_waitrequest)  //                                                     .waitrequest
	);

	mityarm_5csx_dev_board_irq_mapper irq_mapper (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq0_irq)  //    sender.irq
	);

	mityarm_5csx_dev_board_irq_mapper irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (1),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (0),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~hps_0_h2f_reset_reset),         // reset_in0.reset
		.clk            (hps_0_h2f_user0_clock_clk),      //       clk.clk
		.reset_out      (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req      (),                               // (terminated)
		.reset_req_in0  (1'b0),                           // (terminated)
		.reset_in1      (1'b0),                           // (terminated)
		.reset_req_in1  (1'b0),                           // (terminated)
		.reset_in2      (1'b0),                           // (terminated)
		.reset_req_in2  (1'b0),                           // (terminated)
		.reset_in3      (1'b0),                           // (terminated)
		.reset_req_in3  (1'b0),                           // (terminated)
		.reset_in4      (1'b0),                           // (terminated)
		.reset_req_in4  (1'b0),                           // (terminated)
		.reset_in5      (1'b0),                           // (terminated)
		.reset_req_in5  (1'b0),                           // (terminated)
		.reset_in6      (1'b0),                           // (terminated)
		.reset_req_in6  (1'b0),                           // (terminated)
		.reset_in7      (1'b0),                           // (terminated)
		.reset_req_in7  (1'b0),                           // (terminated)
		.reset_in8      (1'b0),                           // (terminated)
		.reset_req_in8  (1'b0),                           // (terminated)
		.reset_in9      (1'b0),                           // (terminated)
		.reset_req_in9  (1'b0),                           // (terminated)
		.reset_in10     (1'b0),                           // (terminated)
		.reset_req_in10 (1'b0),                           // (terminated)
		.reset_in11     (1'b0),                           // (terminated)
		.reset_req_in11 (1'b0),                           // (terminated)
		.reset_in12     (1'b0),                           // (terminated)
		.reset_req_in12 (1'b0),                           // (terminated)
		.reset_in13     (1'b0),                           // (terminated)
		.reset_req_in13 (1'b0),                           // (terminated)
		.reset_in14     (1'b0),                           // (terminated)
		.reset_req_in14 (1'b0),                           // (terminated)
		.reset_in15     (1'b0),                           // (terminated)
		.reset_req_in15 (1'b0)                            // (terminated)
	);

endmodule
